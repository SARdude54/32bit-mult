`timescale 1ps/1ps

module radix4_mult (
    input logic CLK,
    input logic rst_n,
    input logic [32:0] A,
    input logic [32:0] B,
    output logic [32:0] C
);


    
endmodule
